// Generator : SpinalHDL v1.9.3    git head : 029104c77a54c53f1edda327a3bea333f7d65fd9
// Component : Testspinal
// Git hash  : 0508b0a39fa97321c556919db0fe18b82c2b31e4

`timescale 1ns/1ps

module Testspinal (
  input               user_button,
  input               reset_button,
  output reg [5:0]    leds,
  input               xtal_in,
  output              tm_clk,
  inout               tm_dio
);

endmodule
